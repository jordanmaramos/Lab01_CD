library verilog;
use verilog.vl_types.all;
entity LAB01_vlg_check_tst is
    port(
        S1              : in     vl_logic;
        S2              : in     vl_logic;
        S3              : in     vl_logic;
        S4              : in     vl_logic;
        S5              : in     vl_logic;
        S6              : in     vl_logic;
        S7              : in     vl_logic;
        S8              : in     vl_logic;
        S9              : in     vl_logic;
        S10             : in     vl_logic;
        S11             : in     vl_logic;
        S12             : in     vl_logic;
        S13             : in     vl_logic;
        S14             : in     vl_logic;
        S15             : in     vl_logic;
        S16             : in     vl_logic;
        S17             : in     vl_logic;
        S18             : in     vl_logic;
        S19             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end LAB01_vlg_check_tst;
