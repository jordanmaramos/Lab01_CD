library verilog;
use verilog.vl_types.all;
entity LAB01_vlg_check_tst is
    port(
        S1              : in     vl_logic;
        S2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end LAB01_vlg_check_tst;
